LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TECLA IS
PORT(
	CLK,CLR: IN STD_LOGIC;
	F: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	C: INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	DISPLAY: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE A_TECLA OF TECLA IS
CONSTANT TECLA0: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000001";
CONSTANT TECLA1: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001111";
CONSTANT TECLA2: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0010010";
CONSTANT TECLA3: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000110";
CONSTANT TECLA4: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001100";
CONSTANT TECLA5: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100100";
CONSTANT TECLA6: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100000";
CONSTANT TECLA7: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001111";
CONSTANT TECLA8: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000000";
CONSTANT TECLA9: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000100";
CONSTANT TECLANT: STD_LOGIC_VECTOR(6 DOWNTO 0):="0110110";
CONSTANT TECLAG: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001000";
CONSTANT TECLAAST: STD_LOGIC_VECTOR(6 DOWNTO 0):="0110001";
SIGNAL AUX: STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN 
ANILLO: PROCESS(CLK,CLR)
	BEGIN
	IF(CLR='0')THEN
	C<="011";
	ELSIF(CLK'EVENT AND CLK='1')THEN
	C<= TO_STDLOGICVECTOR(TO_BITVECTOR(C) ROR 1);
	END IF;
END PROCESS ANILLO;

DECO: PROCESS(F,C)
BEGIN 
	CASE F&C IS 
	WHEN "1110" & "110" => AUX <= TECLA3;
	WHEN "1101" & "110" => AUX <= TECLA6;
	WHEN "1011" & "110" => AUX <= TECLA9;
	WHEN "0111" & "110" => AUX <= TECLAG;

	WHEN "1110" & "101" => AUX <= TECLA2;
	WHEN "1101" & "101" => AUX <= TECLA5;
	WHEN "1011" & "101" => AUX <= TECLA8;
	WHEN "0111" & "101" => AUX <= TECLA0;

	WHEN "1110" & "011" => AUX <= TECLA1;
	WHEN "1101" & "011" => AUX <= TECLA4;
	WHEN "1011" & "011" => AUX <= TECLA7;
	WHEN "0111" & "011" => AUX <= TECLAAST;
	WHEN OTHERS => AUX<= TECLANT;
END CASE;
END PROCESS DECO;

PROCESS(CLK,CLR,F)
BEGIN
	IF(CLR='0')THEN
		DISPLAY<=TECLANT;
	ELSIF(CLK'EVENT AND CLK='1')THEN
		IF(F="1111")THEN 
			DISPLAY<=DISPLAY;
		ELSE
			DISPLAY<=AUX;
		END IF;
	END IF;
    END PROCESS;
END A_TECLA;


	
	
