LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RC IS 
PORT( CLR,CLK: IN STD_LOGIC;
C,E: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
Q: INOUT STD_LOGIC_VECTOR(2 DOWNTO 0)

);
END ENTITY;

ARCHITECTURE A_RC OF RC IS 
SIGNAL AUX: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL GRAY: STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN 

	conversorGray: process(aux)
	BEGIN 
		gray<=to_stdlogicvector(to_bitvector(aux) xor to_bitvector(aux) srl 1);
	END PROCESS conversorGray;
	
	PROCESS(CLR,CLK,C)
	BEGIN 
	
		IF(CLR='0')THEN
		AUX<="000";
		
		ELSIF(CLK'EVENT AND CLK='1')THEN 
		
			CASE C IS 
				--CARGA DE DATO 
				WHEN "000" => AUX<=E;
				
				--CONTEO ASCENDENTE
				WHEN "001" => AUX<=AUX+1;
				
				--CONTEO DESCENDENTE  
				WHEN "010" => AUX<=AUX-1;
				
				--RETENER
				WHEN "011" => AUX<=AUX;
				
				--CORRIMIENTO A LA DERECHA 
				WHEN "100"=> AUX<=TO_STDLOGICVECTOR(TO_BITVECTOR(AUX) SRL 1);
				
				--CORRIMIENTO A LA IZQUIERDA 
				
				WHEN "101" => AUX<=TO_STDLOGICVECTOR(TO_BITVECTOR(AUX) SLL 1);
				
				--CONTEO ASCENDENTE GRAY 
				WHEN "110" => AUX<=AUX+1;
				
				--CONTEO DESCENDENTE GRAY 
				WHEN OTHERS => AUX<=AUX-1;
				
			END CASE;
		END IF
	END PROCESS;
	
	PROCESS(C,GRAY,AUX)
	BEGIN 
		IF(C="110" OR C="111")THEN 
			Q<=GRAY;
		ELSE 
			Q<=AUX;
		END IF;
	END PROCESS;
END A_RC;
			