LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ContadorD IS 
PORT(CLK, CLR, C: IN STD_LOGIC;
     Q: INOUT STD_LOGIC_VECTOR (2 DOWNTO 0));
END ENTITY;

ARCHITECTURE A_ContadorD OF ContadorD IS 
SIGNAL D: STD_LOGIC_VECTOR (2 DOWNTO 0);
BEGIN
     PROCESS(C, Q)
	 BEGIN
	      D(2) <= (C AND Q(2)) OR (Q(2) AND NOT Q(1)) OR (Q(2)AND NOT Q(0)) OR (NOT C AND NOT Q(2) AND Q(1) AND Q(0));
          D(1) <= (Q(1) AND NOT Q(0)) OR (C AND Q(1)) OR (NOT C AND NOT Q(1) AND Q(0));
		  D(0) <= C XNOR Q(0);
	 END PROCESS;

     PROCESS(CLK, CLR)
	 BEGIN
	      IF (CLR = '0')THEN
		  Q <= "000";
	 ELSIF(CLK'EVENT AND CLK='1')THEN
	      Q <= D;
	 END IF;
	END PROCESS;
 END A_ContadorD;