LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONDEC IS
	PORT(CLK, CLR : IN STD_LOGIC;
			C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			E: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DISPLAY: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);

ATTRIBUTE PIN_NUMBERS OF CONDEC : ENTITY IS
"CLK:1 CLR:2 C(1):3 C(0):4 E(3):5 E(2):6 E(1):7 E(0):8";
END ENTITY;
ARCHITECTURE A_CONDEC OF CONDEC IS
	CONSTANT DIG0 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000001";
	CONSTANT DIG1 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001111";
	CONSTANT DIG2 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0010010";  
	CONSTANT DIG3 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000110";
	CONSTANT DIG4 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001100";
	CONSTANT DIG5 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100100";
	CONSTANT DIG6 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100000";
	CONSTANT DIG7 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001111";
	CONSTANT DIG8 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000000";
	CONSTANT DIG9 : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000100";
BEGIN
	PROCESS(CLR, CLK,C, DISPLAY)
	BEGIN
		IF(CLR='0') THEN
			DISPLAY <= DIG0;
		ELSIF (CLK'EVENT AND CLK='1') THEN
			CASE C IS
				WHEN "00"=> --Contador ascendente
					CASE DISPLAY IS
						WHEN DIG0 => DISPLAY <= DIG1;
						WHEN DIG1 => DISPLAY <= DIG2;
						WHEN DIG2 => DISPLAY <= DIG3;
						WHEN DIG3 => DISPLAY <= DIG4;
						WHEN DIG4 => DISPLAY <= DIG5;
						WHEN DIG5 => DISPLAY <= DIG6;
						WHEN DIG6 => DISPLAY <= DIG7;
						WHEN DIG7 => DISPLAY <= DIG8;
						WHEN DIG8 => DISPLAY <= DIG9;
						WHEN OTHERS => DISPLAY <= DIG0;
					END CASE;
				WHEN "01"=> --Contador Descendente
					CASE DISPLAY IS
					    WHEN DIG0 => DISPLAY <= DIG9;
						WHEN DIG9 => DISPLAY <= DIG8;
						WHEN DIG8 => DISPLAY <= DIG7;
						WHEN DIG7 => DISPLAY <= DIG6;
						WHEN DIG6 => DISPLAY <= DIG5;
						WHEN DIG5 => DISPLAY <= DIG4;
						WHEN DIG4 => DISPLAY <= DIG3;
						WHEN DIG3 => DISPLAY <= DIG2;
						WHEN DIG2 => DISPLAY <= DIG1;	
						WHEN OTHERS => DISPLAY <= DIG0;
					END CASE;
				WHEN "10"=>DISPLAY<=DISPLAY; --Retener Dato
					
				WHEN OTHERS => 
					CASE E IS
						WHEN "0000" => DISPLAY <= DIG0;
						WHEN "0001" => DISPLAY <= DIG1;
						WHEN "0010" => DISPLAY <= DIG2;
						WHEN "0011" => DISPLAY <= DIG3;
						WHEN "0100" => DISPLAY <= DIG4;
						WHEN "0101" => DISPLAY <= DIG5;
						WHEN "0110" => DISPLAY <= DIG6;
						WHEN "0111" => DISPLAY <= DIG7;
						WHEN "1000" => DISPLAY <= DIG8;
						WHEN OTHERS => DISPLAY <= DIG9;
					END CASE;
			END CASE;
		END IF;
	END PROCESS;
END A_CONDEC;
