module entdeco ( 
	entry,
	display
	) ;

input [1:0] entry;
inout [6:0] display;
