LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONTADOR_8B IS
	PORT
	(
		CLK,CLR: IN STD_LOGIC;
		CONTROL: IN STD_LOGIC;
		Q: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)	-- Se puede ocupar el 2 1 0
	);

END ENTITY;


ARCHITECTURE A_CONT OF CONTADOR_8B IS
SIGNAL J_Y_K: STD_LOGIC_VECTOR(7 DOWNTO 0);	--AQU� IRAN LAS ENTRADAS J Y K DEL FLIP-FLOP EN UNA SIGNAL 
--LA SIGANLS CAMBIAN DE VALOR HASTA QUE LAS TERMINA DE USAR UN PROCESO
BEGIN 
	
	-- LOS PROCESS INDICAN UN ORDEN, SER�AN COMO BLOQUES DE C�DIGO EN C, JAVA, ETC.
	COMP_AND:PROCESS(CONTROL,Q)	-- LOS ARGUMENTOS DE LA LISTA SENSITIVA O EL PROCESS SON OPCIONALES
	BEGIN
		J_Y_K(7)<=(NOT CONTROL)AND(Q(6))AND(Q(5))AND(Q(4))AND(Q(3))AND(Q(2))AND(Q(1))AND(Q(0));
		J_Y_K(6)<=(NOT CONTROL)AND(Q(5))AND(Q(4))AND(Q(3))AND(Q(2))AND(Q(1))AND(Q(0));
		J_Y_K(5)<=(NOT CONTROL)AND(Q(4))AND(Q(3))AND(Q(2))AND(Q(1))AND(Q(0));
		J_Y_K(4)<=(NOT CONTROL)AND(Q(3))AND(Q(2))AND(Q(1))AND(Q(0));
		J_Y_K(3)<=(NOT CONTROL)AND(Q(2))AND(Q(1))AND(Q(0));
		J_Y_K(2)<=(NOT CONTROL)AND(Q(1))AND(Q(0));
		J_Y_K(1)<=(NOT CONTROL)AND(Q(0));
		J_Y_K(0)<=(NOT CONTROL);
	END PROCESS COMP_AND;
	
	-- IMPLEMENTANDO EL FLIP-FLOP JK
	FF_JK:process(CLR,CLK,Q,J_Y_K)
	BEGIN
		IF(CLR='0')THEN
			Q<="00000000";
		ELSIF(CLK'EVENT AND CLK='1')THEN
			Q<=(J_Y_K AND NOT Q)OR(NOT J_Y_K AND Q);
		END IF;
	end PROCESS FF_JK;

END A_CONT;